library ieee;
use ieee.std_logic_1164.all;

entity Datapath is
	port (
		return_all : in std_logic;
	)