LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

-- MEMÓRIA EEPROM
ENTITY EEPROM IS
	GENERIC (
		ADDR_LENGHT : NATURAL := 4;
		R_LENGHT : NATURAL := 8;
		NUM_OF_REGS : NATURAL := 16
	);
	PORT (
		clk : IN STD_LOGIC;
		wr : IN STD_LOGIC;
		addr : IN STD_LOGIC_VECTOR (ADDR_LENGHT - 1 DOWNTO 0);
		datain : IN STD_LOGIC_VECTOR (R_LENGHT - 1 DOWNTO 0);
		dataout : OUT STD_LOGIC_VECTOR (R_LENGHT - 1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE ROM_REGISTER OF EEPROM IS
	TYPE rom_reg IS ARRAY (0 TO NUM_OF_REGS - 1) OF
	STD_LOGIC_VECTOR (R_LENGHT - 1 DOWNTO 0);
	SIGNAL rom_s : rom_reg;

	begin
		process(clk)
		variable loc : integer;
		begin
			if (rising_edge(clk)) then
				loc := to_integer(unsigned(addr));
				if (wr = '1') then
					rom_s(loc) <= datain;
				end if;
				dataout <= ram_s(loc);
			end if;
		end process;
end architecture ROM_REGISTER;
